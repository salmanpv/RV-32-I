package Types;

typedef Bit#(32) Word;
typedef Bit#(5)  RegIdx;
typedef Bit#(7)  Opcode;
typedef Bit#(3)  Funct3;
typedef Bit#(7)  Funct7;
typedef Bit#(1)  Bit1;

endpackage

